`ifndef _AD9958_VARS_VH_

`define _AD9958_VARS_VH_

`define IOMODE_2_WIRE 2'b00
`define IOMODE_3_WIRE 2'b01
`define IOMODE_2_BIT 2'b10
`define IOMODE_4_BIT 2'b11

`define DAC_FSCALE_FULL 2'b11
`define DAC_FSCALE_HALF 2'b01
`define DAC_FSCALE_QUARTER 2'b10
`define DAC_FSCALE_EIGHTH 2'b00

`endif
