/*
 * Registers accessed in this project is listed here.
 */

`ifndef _AD9958_ADDRESS_VH_

`define _AD9958_ADDRESS_VH_

`define ADDR_CSR 8'h00
`define ADDR_FR1 8'h01
`define ADDR_FR2 8'h02
`define ADDR_CFR 8'h03
`define ADDR_CFTW0 8'h04
`define ADDR_ACR 8'h06

`endif
